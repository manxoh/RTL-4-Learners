module axis_pipe #(AXIS_WIDTH = 32)
                                  (input clk,
                                   input reset,
                                   input s_axis_tvalid,
                                   input [AXIS_WIDTH-1:0] s_axis_tdata,
                                   output s_axis_tready,
                                   output m_axis_tvalid,
                                   output [AXIS_WIDTH-1:0] m_axis_tdata,
                                   input m_axis_tready);

   //internal signals

   //modify data

   //outputs

endmodule
