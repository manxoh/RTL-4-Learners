module axis_sink #(AXIS_WIDTH = 32)
                                  (input clk,
                                   input reset,
                                   input s_axis_tvalid,
                                   input [AXIS_WIDTH-1:0] s_axis_tdata,
                                   output s_axis_tready,
                                   output valid,
                                   output [AXIS_WIDTH-1:0] data_out);

   //internal signals

   //modify data

   //outputs

endmodule
